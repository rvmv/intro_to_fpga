
module board_terasic
(
    input         CLK,
    input  [ 9:0] SW,
    input  [ 1:0] KEY,
    output [ 9:0] LED,
    output [ 7:0] HEX0,
    output [ 7:0] HEX1,
    output [ 7:0] HEX2,
    output [ 7:0] HEX3,
    output [ 7:0] HEX4,
    output [ 7:0] HEX5 
);

//switch_to_led sw_to_led (.SW(SW), .LEDR(LED));

//mux_2_to_1_simple mux (.SW(SW), .LEDR(LED));

//mux_2_to_1_procedural mux_procedural (.SW(SW), .LEDR(LED));

knight_rider kr (.CLOCK_50(CLK), .LEDR(LED), .SW(SW));

endmodule